
Installation
------------
 
Detta Arkiv inneh�ller det Svenska Spr�kst�det (NLS) f�r
XWorkplace. Det f�ruts�tter att en installerad XWP Version 0.9.20
finns p� systemet.
 
P� den sista sidan "System Konfiguration" kan man best�mma, om
WarpIN skall skapa WPS-Objekt, f�r XWorkplace och den Svenska 
Spr�kversionen. Aktivera Optionen "Skapa WPS objekt". Beakta ocks�
anm�rkningen under Punkt 1 hos "K�nda Problem". Det g�r ocks�
att vid ett senare tillf�lle skapa Svenska objekt och menyer
genom att k�ra de bifogade REXX-Scripten "instl046.cmd", "crobj06.cmd"
och "sound046.cmd" i underkatalogen install hos XWorkplace.
 
N�r paketet har installerats med WarpIN, m�ste det Svenska spr�ket
aktiveras p� f�ljande s�tt:
 
1. �ppna Objektet "XWorkplace Setup".
2. V�lj fliken med "XWorkplace Status".
3. V�lj i rullningslisten under "National Language Support" 
   alternativet "SV Svenska -- xfldr046.dll".
4. Bekr�fta �ndringen i Dialogen, och st�ng Notboken. N�sta g�ng den
   �ppnas �r spr�ket �ndrat.
 
 
K�nda Problem och Inskr�nkningar
--------------------------------
 
1. Genom uppst�llningen hos Konfigurations-Ordningen hos de
   Svenska Objektrubrikerna kan de tidigare gjorda personliga
   inst�llningarna och menyalternativen f�rloras.

2. N�r Spr�kversioner �ndras via Objektet "XWorkplace-Setup", 
   kan det f�rekomma att XCenter inte f�ljer med och �ndras till
   r�tt Spr�k. Detta kan l�sas genom att st�nga av och starta om 
   XCenter en g�ng.
 
 
Kontakter
---------
 
Har n�gon problem med det Engelska spr�ket eller om ni hittar n�got
fel i �vers�ttningen, skicka ett E-mail till �vers�ttaren
Bj�rn S�derstr�m p� adress: bjorso@os2ug.se

F�r �vriga �renden om fel i sj�lva XWorkplace etc. h�nvisas till de
speciella mailinglistor som finns f�r XWorkplace. L�s i den bifogade 
Anv�ndarguiden om adresser till listorna. XWorkplace �r en produkt som
utvecklas snabbt och d�rf�r kan man inte vara helt s�ker p� att den 
fungerar helt perfekt med alla kombinationer av h�rdvara, spr�k, revl�gen p� 
operativsystemet m.m. I de allra flesta fall fungerar den mycket bra
och det finns gott om tips i dokumentationen om problem skulle uppst�.

Anm�rkning: 
         Det Svenska Spr�kst�det f�r XWorkplace har i m�jligaste m�n
	 f�ljt standard hos OS/2 och eCS. F�r �mnen d�r en �vers�ttning
	 inte skulle f�rb�ttra en Svensk version har orginalengelskan 
	 beh�llits. Eftersom den etablerade terminologin f�r data och datorer
	 �r Engelska skulle en f�rsvenskning av tekniska termer troligtvis vara
	 till det s�mre f�r de flesta anv�ndare. 
 
Nerladdning
--------
 
Aktuell Version av Spr�kpaketet kan h�mtas med f�ljande URL l�nk:
 
http://www.os2ug.se/zippar/xwp-0-9-20_nls_sv.exe
 
K�llkoden f�r spr�ket finns tillg�nglig p� XWorkplace-CVS-Arkiv hos
Netlabs (Under katalogen 046). H�nvisning f�r hur dessa Arkiv nyttjas
finns under adressen http://www.xworkplace.org/cvs.html.
 
Datum: 12/11/2002
